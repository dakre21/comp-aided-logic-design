`timescale 1ns / 1ns

// HLS has generated this HDL code with the hlsyn executable
// Author: David Akre

module HLSM (Clk, Rst, Start, Done);
    input Clk, Rst, Start;
    output reg Done;
     reg [31:0] a, b, c, d, e, f, g, h, sa;
      reg [31:0] avg;
      reg [31:0] t1, t2, t3, t4, t5, t6, t7, t7div2, t7div4;


// Initial Wait State S0 of the HLSM
    always @(posedge Clk, ~Start) begin
    // Do nothing
    end

// C to HLSM states below based on FDS scheduling
    always @(posedge Clk, a, b, c, t1, Start) begin
        t1 = a + b;
        t2 = t1 + c ;
    end

    always @(posedge Clk, d, t2) begin
        t3 = t2 + d ;
    end

    always @(posedge Clk, e, t3) begin
        t4 = t3 + e ;
    end

    always @(posedge Clk, f, t4) begin
        t5 = t4 + f ;
    end

    always @(posedge Clk, g, t5) begin
        t6 = t5 + g ;
    end

    always @(posedge Clk, h, t6) begin
        t7 = t6 + h ;
    end

    always @(posedge Clk, a, sa) begin
        t7div2 = t7 >> sa;
    end

    always @(posedge Clk, a, sa, t7div2) begin
        t7div4 = t7div2 >> sa ;
    end

    always @(posedge Clk, d, sa, t7, t7div4) begin
        avg = t7div4 >> sa;
    end

// Final State to conclude the HLSM by setting Done to logic level high (i.e. 1)
    always @(posedge Clk,  avg ) begin
        Done = 1;
    end


endmodule
